module top_module(
    input [1023:0] in,
    input [7:0] sel,
    output [3:0] out );
    assign out = in[sel*4+3 -: 4];
endmodule
//
//答案
//
//assign out = {in[sel*4+3], in[sel*4+2], in[sel*4+1], in[sel*4+0]};
    // We can't part-select multiple bits without an error, but we can select one bit at a time,
    // four times, then concatenate them together.
    //
    // Alternatively, "indexed vector part select" works better, but has an unfamiliar syntax:
    // assign out = in[sel*4 +: 4];        // Select starting at index "sel*4", then select a total width of 4 bits with increasing (+:) index number.
    // assign out = in[sel*4+3 -: 4];    // Select starting at index "sel*4+3", then select a total width of 4 bits with decreasing (-:) index number.
    // Note: The width (4 in this case) must be constant.